// REQUIREMENTS:
// 	This module turns a 2D array into 8 outputs for the sr_ctrl
// 	Handles an LED reset, doesnt send anything for 50us
// 